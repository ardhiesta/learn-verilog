//dataflow and gate with two inputs
module and2 (x1, x2, z1);

input x1, x2;
output z1;

wire x1, x2;
wire z1;

assign z1 = x1 & x2;

endmodule
